module PC_Adder (
    input [63:0]a,b,
    output [63:0]c
);

    assign c = a + b;
    
endmodule